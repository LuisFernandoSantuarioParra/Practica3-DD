LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
LIBRARY LATTICE;
USE LATTICE.ALL;
use ieee. std_logic_arith.all;
use ieee. std_logic_unsigned.all;

ENTITY FFPORTS IS

	PORT(
			
		CLK,CLR,J,K,S,R,D,T:IN STD_LOGIC;		
		SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		DISPLAY: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
	
END FFPORTS;
ARCHITECTURE FFPROGRAMS OF FFPORTS IS

SIGNAL QD,QJK,QT,QRS,Q: STD_LOGIC;
BEGIN
		PFFD:PROCESS(CLK,CLR)
		BEGIN
			IF(CLR='1')THEN
				QD<='0';
			ELSIF(CLK'EVENT AND CLK='1') THEN
				QD<=D;
			END IF;
		END PROCESS PFFD;
		
		
		PFFJK:PROCESS(CLK,CLR)
		BEGIN
			IF(CLR='1')THEN
				QJK<='0';
			ELSIF(CLK'EVENT AND CLK='1') THEN
				QJK<=(NOT K AND QJK) OR (J AND NOT QJK);
			END IF;
		END PROCESS PFFJK;
		
		
		PFFRS:PROCESS(CLK)
		BEGIN
		
			IF(CLK'EVENT AND CLK='1') THEN
				
				IF(S='0' AND R='1')THEN
					QRS<='0';
				ELSIF(S='1' AND R='0')THEN
					QRS<='1';
				ELSIF(S='0' AND R='0')THEN
					QRS<=QRS;
				END IF;
				
			END IF;
		END PROCESS PFFRS;
		
		
		PFFT:PROCESS(CLK)
		BEGIN
			IF(CLK'EVENT AND CLK='1') THEN
				IF T='0' THEN
					QT <= QT;
					ELSIF T='1' THEN
					QT <= not (QT);
					END IF;
			END IF;
		END PROCESS PFFT;
		
		
	WITH SEL SELECT
		Q <= QD  WHEN "00" , 
		    QJK  WHEN "01" ,
		    QT   WHEN "10" ,
		    QRS  WHEN OTHERS;

DISPLAY <="0000001" WHEN (Q='0')ELSE
			"1001111";


END FFPROGRAMS;